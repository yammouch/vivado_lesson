module sim_top;

initial begin
  $display(`SCENARIO_NAME);
end

`include `SCENARIO_NAME

endmodule
