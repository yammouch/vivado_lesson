module sub (
 input  di,
 output do );

assign do = !di;

endmodule
