architecture sim2 of sim_top is
begin
  process
  begin
    report "sim2";
    wait;
  end process;
end sim2;
