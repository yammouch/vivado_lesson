entity sim_top is
end entity;
