initial begin
  $display("s02");
end
