architecture sim1 of sim_top is
begin
  process
  begin
    report "sim1";
    wait;
  end process;
end sim1;
