initial begin
  $display("s01");
end
